
`ifndef AHB_AGENT_PKG_SV
`define AHB_AGENT_PKG_SV

`include "ahb_if.sv"

package agent_pkg;


  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  `include "../src/agent/transaction.sv"
  `include "../src/agent/seq_item.sv"
  `include "../src/agent/sequence.sv"
  `include "../src/agent/sequencer.sv"
  `include "../src/agent/driver.sv"
  `include "../src/agent/monitor.sv"
  `include "../src/agent/agent_config.sv"
  `include "../src/agent/agent.sv"
  `include "../src/agent/env.sv"
  `include "../src/agent/test.sv"
  
endpackage: agent_pkg;
  
`endif