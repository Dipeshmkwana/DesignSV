
class apb3_ms_testcase_config;
  
  function new();
  endfunction
endclass
