package apb3_ms_pkg;
`include "../src/apb3_ms_agent/apb3_ms_txn.sv"
`include "../src/apb3_ms_agent/apb3_m_generator.sv"
`include "../src/apb3_ms_agent/apb3_ms_functional_coverage.sv"
`include "../src/apb3_ms_agent/apb3_m_driver.sv"
`include "../src/apb3_ms_agent/apb3_m_monitor.sv"
`include "../src/apb3_ms_agent/apb3_m_agent.sv"
`include "../src/apb3_ms_agent/apb3_s_generator.sv"
`include "../src/apb3_ms_agent/apb3_s_driver.sv"
`include "../src/apb3_ms_agent/apb3_s_monitor.sv"
`include "../src/apb3_ms_agent/apb3_s_agent.sv"
`include "../src/apb3_ms_agent/apb3_ms_env.sv"
`include "../src/apb3_ms_agent/apb3_ms_testcase.sv"
`include "../src/apb3_ms_agent/apb3_ms_interface.sv"
endpackage


