//----------------
// ABP Design
//----------------
//  Module: apb3
//
module apb3
  /*  package imports  */
  #(
    WIDTH
  )(
    PCLK,
    PRESETn,
    PSLVERR,
    PREADY,
    
  );

  
endmodule: apb3
