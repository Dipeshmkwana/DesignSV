/* -.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-. 
* File Name     : env_cofig.sv
* File Directory: env
* Description   : 
* Author        : Dipesh Makwana 
* Creation Date : 28-05-2019
* Last Modified : Tuesday 28 May 2019 12:12:53 PM IST
* Organization  : Eitra 
* Copyright (c) 2019 Eitra. All rights reserved.
* -.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-.-. */ 
class apb3_ms_env_config_c;

  function new();
    
  endfunction

endclass
