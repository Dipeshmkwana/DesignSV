class apb3_ms_env_config_c;

  function new();
    
  endfunction

endclass