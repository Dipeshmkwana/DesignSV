package base_pkg;


  import uvm_pkg::*;
  `include "uvm_macros.svh"
  
  // `include "base_transaction.sv"
  // `include "base_seq_1.sv"
  // `include "base_sequence.sv"
  // `include "base_sequencer.sv"
  // `include "base_driver.sv"
  // `include "base_monitor.sv"
  // `include "base_agent_config.sv"
  // `include "base_agent.sv"
  // `include "base_env.sv"
  // `include "base_test.sv"
  
  endpackage: base_pkg;