package ahb_env_pkg;

  `include "ahb_env.sv"
  `include "ahb_if.sv"
  
  
endpackage: ahb_env_pkg;