

// suppose it is for APB vip

module top_tb;
  //import uvm pkg

  //declaration
  bit PCLK;
  bit PRESETn;
  wire PSLVERR;
  wire PREADY;
  wire PWRITE;
  wire PENABLE;
  wire PSELx;
  wire[31:0] PADDR;
  wire[31:0] PWDATA;
  wire[31:0] PRDATA;
  wire PSTRB;
  wire PPROT;

  //interface declaration
  

  // environment instance 

  // DUT instance 

  //Clock init

  //UVM Start up

  //Dump waves

endmodule : top_tb

