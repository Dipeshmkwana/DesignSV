package ahb_vip_pkg;

  `include "ahb_agent.sv"
  `include "ahb_scoreboard"
  `include "ahb_monitor"
  
endpackage: ahb_vip_pkg;