// copyright 2014 definitely_launch inc.
// Description	:
// creation date: 
// modified date: 
// Authored by  : Vinod Sureshkumar Ailsinghani
// Fie Name	: 
// version	: 1.0

package skeleton_env;


import uvm_pkg::*;
`include "uvm_macros.svh"

/*`include "asic_jan2018_transaction.sv"
`include "asic_jan2018_seq_1.sv"
`include "asic_jan2018_sequencer.sv"
`include "asic_jan2018_driver.sv"
`include "asic_jan2018_monitor.sv"
`include "asic_jan2018_agent_config.sv"
`include "asic_jan2018_agent.sv"
`include "asic_jan2018_env.sv"
`include "asic_jan2018_test.sv"
*/

endpackage
