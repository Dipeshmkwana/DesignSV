 // Sequence item contains the data 
  class base_seq_item extends uvm_sequence_item;
    
  endclass: base_pkg